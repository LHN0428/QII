library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SHFTB IS 

PORT (CLK,LOAD,SR:IN STD_LOGIC ;
		 DIN :IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
		 QB :OUT STD_LOGIC ;
		 DOUT :OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);
END SHFTB;

ARCHITECTURE behav OF SHFTB IS 
SIGNAL REG8 :STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
PROCESS(CLK,LOAD)
BEGIN
    IF LOAD = '1' THEN 
        REG8 <= DIN ;
		  ELSE IF CLK'EVENT AND CLK = '1' THEN
		  REG8(6 DOWNTO 0 )<= REG8(7 DOWNTO 1) ;
    	 END IF ;
    END IF ;
		  END PROCESS ;
		  QB <=REG8(0) ;
		  DOUT <= SR & REG8(7 DOWNTO 1) ;
		  END behav;