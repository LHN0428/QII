library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY cnt9 IS
port (CLK,RST,EN:IN STD_LOGIC;
			COUT : OUT STD_LOGIC
	   );

END cnt9;
			
ARCHITECTURE behav OF cnt9 IS
BEGIN 
	PROCESS (CLK,RST,EN)
	VARIABLE Q:STD_LOGIC_VECTOR(3 DOWNTO 0);
	BEGIN
	
	IF RST = '0'  THEN Q:="0001" ;
	ELSIF CLK'EVENT AND CLK='1' THEN
			IF EN='0' THEN 
			IF Q<"1010" THEN Q:=Q+1 ;
			ELSE Q:="0001" ;
			END IF ;
		END IF;
	 END IF ;
 
 IF Q="1010" THEN COUT <='1';
 ELSE COUT<='0' ;
 END IF ;
 
 END PROCESS;
 END behav ;
 

			

