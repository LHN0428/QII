library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY dffen IS

PORT(EN:IN STD_LOGIC;
      D: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		Q: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	 );
END dffen ;

ARCHITECTURE behav OF dffen IS
BEGIN
PROCESS(D,EN)
BEGIN
IF EN='0' THEN Q <= (OTHERS =>'0');
ELSE Q<=D;
END IF ;
END PROCESS ;
END behav ;