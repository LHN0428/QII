library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SHFTA IS 

PORT (CLK,CLR,SR:IN STD_LOGIC;
		DIN : IN STD_LOGIC_VECTOR (7 DOWNTO 0) ;
		QB :  OUT STD_LOGIC ;
		DOUT : OuT STD_LOGIC_VECTOR (7 DOWNTO 0));
END SHFTA ;

ARCHITECTURE behav OF SHFTA IS
 
SIGNAL REG8:STD_LOGIC_VECTOR (7 DOWNTO 0);
SIGNAL Q:STD_LOGIC ;

BEGIN
PROCESS (CLK ,CLR)
BEGIN 
	IF CLR = '1' THEN 
	REG8 <= (OTHERS=>'0') ;  
	Q <= '0';
	ELSIF CLK'EVENT AND CLK ='1' THEN
	REG8 <= DIN;
	Q <=SR ;
	END IF ;
	DOUT <= Q & REG8(7 DOWNTO 1) ;    
	END PROCESS ;
	QB <= REG8(0) ;
	END behav ;
	
	